// This file is public domain, it can be freely copied without restrictions.
// SPDX-License-Identifier: CC0-1.0

module dut ( 
  input                       aclk,
  input                       arstn
);


endmodule
